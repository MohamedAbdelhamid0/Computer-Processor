--
--	Package File Template
--
--	Purpose: This package defines supplemental types, subtypes, 
--		 constants, and functions 
--
--   To use any of the example code shown below, uncomment the lines and modify as necessary
--

library IEEE;
use IEEE.STD_LOGIC_1164.all;
USE IEEE.NUMERIC_STD.ALL;


package decoderpack is

component decoder is
 Port ( s : in  STD_LOGIC_VECTOR (4 downto 0);
			  l0: out STD_LOGIC;
			  l1: out STD_LOGIC;
			  l2: out STD_LOGIC;
			  l3: out STD_LOGIC;
			  l4: out STD_LOGIC;
			  l5: out STD_LOGIC;
			  l6: out STD_LOGIC;
			  l7: out STD_LOGIC;
			  l8: out STD_LOGIC;
			  l9: out STD_LOGIC;
			  l10: out STD_LOGIC;
			  l11: out STD_LOGIC;
			  l12: out STD_LOGIC;
			  l13: out STD_LOGIC;
			  l14: out STD_LOGIC;
			  l15: out STD_LOGIC;
			  l16: out STD_LOGIC;
			  l17: out STD_LOGIC;
			  l18: out STD_LOGIC;
			  l19: out STD_LOGIC;
			  l20: out STD_LOGIC;
			  l21: out STD_LOGIC;
			  l22: out STD_LOGIC;
			  l23: out STD_LOGIC;
			  l24: out STD_LOGIC;
			  l25: out STD_LOGIC;
			  l26: out STD_LOGIC;
			  l27: out STD_LOGIC;
			  l28: out STD_LOGIC;
			  l29: out STD_LOGIC;
			  l30: out STD_LOGIC;
			  l31: out STD_LOGIC );	  

end component;


end decoderpack;

